module DeNoiser();

endmodule